


module mul(
    input wire 
    input wire 
    input wire
    input wire
);

endmodule